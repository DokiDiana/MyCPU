module FORWARD(
    input IDEX_rs1,
    input IDEX_rs2,
    input EXMEM_RegWrite,
    input EXMEM_rd,
    input MEMWB_RegWrite,
    input MEMWB_rd,
    output F1, F2,
);